B8201073B0201073
4201418141014081
4401438143014281
4601458145014481
4801478147014681
4A01498149014881
4C014B814B014A81
4E014D814D014C81
53374F814F014E81
1073555303135555
8193000031977C03
0113000031178EE1
0513000025170E61
8593000025970DE5
202300B577630D65
FEB56DE305110005
2029458145012091
000000000000A001
FFFE0E1300010E37
408E8E9380001EB7
800015B701CEA023
0005A28340058593
4045051380001537
005520230102D293
C4221141FE0002E3
041300000417C04A
091300000917F364
C60640890933F2E9
096340295913C226
0485401C44810009
FE991CE397820411
F084041300000417
F009091300000917
4029591340890933
401C448100090963
1CE3978204110485
4492442240B2FE99
0000808201414902
0000000000000000
